package async_fifo_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "sv_fifo_sequence_item.svh"
    `include "sv_fifo_sequence.svh"

    `include "sv_fifo_monitor.svh"
    `include "sv_fifo_driver.svh"
    `include "sv_fifo_scoreboard.svh"
    `include "sv_fifo_sequencer.svh"
    `include "sv_fifo_virtual_sequencer.svh"
    `include "sv_fifo_agent.svh"
    `include "sv_fifo_env.svh"

    `include "sv_case_sequence.svh"

    `include "sv_base_test.svh"
    `include "sv_case_test.svh"

endpackage